/////////////////////////////////////////////////////
// Module interface
/////////////////////////////////////////////////////

module lm32_dp_ram(
	// ----- Inputs -----
	clk_i,
	rst_i,
	we_i,
	waddr_i,
	wdata_i,
	raddr_i,
	// ----- Outputs -----
	rdata_o
);

/////////////////////////////////////////////////////
// Parameters
/////////////////////////////////////////////////////

parameter data_width = 1;               // Width of the data ports
parameter addr_width = 1;               // Width of the address ports

/////////////////////////////////////////////////////
// Inputs
/////////////////////////////////////////////////////

input clk_i;
input rst_i;
input we_i;
input [addr_width-1:0] waddr_i;
input [data_width-1:0] wdata_i;
input [addr_width-1:0] raddr_i;

/////////////////////////////////////////////////////
// Outputs
/////////////////////////////////////////////////////

output [data_width-1:0] rdata_o;

/////////////////////////////////////////////////////
// Internal nets and registers
/////////////////////////////////////////////////////

reg [data_width-1:0] mem[(1<<addr_width)-1:0];
reg [addr_width-1:0] raddr_r;

/////////////////////////////////////////////////////
// Combinational logic
/////////////////////////////////////////////////////

assign rdata_o = mem[raddr_r];

/////////////////////////////////////////////////////
// Sequential logic
/////////////////////////////////////////////////////

integer i;

initial
begin
	for (i = addr_depth-1 ; i >= 0 ; i = i-1)
	begin
		ram[i] <= {data_width{1'b0}};
	end
end

always @(posedge clk_i)
begin
	if (we_i)
		mem[waddr_i] <= wdata_i;
	raddr_r <= raddr_i;
end

endmodule

